VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
	LAYER LEF58_BACKSIDE STRING ;
	LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

LAYER OVERLAP
	TYPE OVERLAP ;
END OVERLAP

LAYER MB
	TYPE ROUTING ;
	PROPERTY LEF58_BACKSIDE "BACKSIDE ; " ;
	DIRECTION HORIZONTAL ;
	PITCH   300 ;
	WIDTH   60 ;
	SPACING 180  ;
END MB

LAYER TSV1
	TYPE CUT ;
	PROPERTY LEF58_TYPE "TYPE TSV ; " ;
END TSV1

LAYER METAL1
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 0.3 ;
	SPACING 0.3 ;
	PITCH 0.6 ;
	MINIMUMCUT 2 WIDTH 1.5 FROMABOVE ;
END METAL1

LAYER VIA12
	TYPE CUT ;
	SPACING 0.4 ;
END VIA12

LAYER METAL2
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 0.3 ;
	SPACING 0.3 ;
	PITCH 0.6 ;
	MINIMUMCUT 2 WIDTH 1.5 ;
END METAL2

LAYER VIA23
	TYPE CUT ;
	SPACING 0.4 ;
END VIA23

LAYER METAL3
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 0.3 ;
	SPACING 0.3 ;
	PITCH 0.6 ;
	MINIMUMCUT 2 WIDTH 1.5 ;
END METAL3

LAYER VIA34
	TYPE CUT ;
	SPACING 0.4 ;
END VIA34

LAYER METAL4
	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	WIDTH 0.3 ;
	SPACING 0.3 ;
	PITCH 0.6 ;
	MINIMUMCUT 2 WIDTH 1.5 FROMBELOW ;
END METAL4

LAYER VIA45
	TYPE CUT ;
	SPACING 1.8 ;
END VIA45

LAYER RDL
	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	WIDTH 2.8 ;
	SPACING 1.8 ;
	PITCH 5.4 ;
	MAXWIDTH 30 ;
END RDL

VIA VIA_TSV
	LAYER MB ;
		RECT -25 -25 25 25 ;
	LAYER TSV1 ;
		RECT -6.5 -6.5 6.5 6.5 ;
	LAYER METAL1 ;
		RECT -6.5 -6.5 6.5 6.5 ;
END VIA_TSV

VIA VIA12_1 DEFAULT
	LAYER METAL1 ;
		RECT -0.3 -0.3 0.3 0.3 ;
	LAYER VIA12 ;
		RECT -0.15 -0.15 0.15 0.15 ;
	LAYER METAL2 ;
		RECT -0.3 -0.3 0.3 0.3 ;
END VIA12_1

VIA VIA12_2H DEFAULT
	LAYER METAL1 ;
		RECT -0.75 -0.3 0.75 0.3 ;
	LAYER VIA12 ;
		RECT -0.6 -0.15 -0.3 0.15 ;
		RECT 0.3 -0.15 0.6 0.15 ;
	LAYER METAL2 ;
		RECT -0.75 -0.3 0.75 0.3 ;
END VIA12_2H

VIA VIA12_2V DEFAULT
	LAYER METAL1 ;
		RECT -0.3 -0.75 0.3 0.75 ;
	LAYER VIA12 ;
		RECT -0.15 -0.6 0.15 -0.3 ;
		RECT -0.15 0.3 0.15 0.6 ;
	LAYER METAL2 ;
		RECT -0.3 -0.75 0.3 0.75 ;
END VIA12_2V

VIA VIA12_4 DEFAULT
	LAYER METAL1 ;
		RECT -0.75 -0.75 0.75 0.75 ;
	LAYER VIA12 ;
		RECT -0.6 -0.6 -0.3 -0.3 ;
		RECT -0.6 0.3 -0.3 0.6 ;
		RECT 0.3 0.3 0.6 0.6 ;
		RECT 0.3 -0.6 0.6 -0.3 ;
	LAYER METAL2 ;
		RECT -0.75 -0.75 0.75 0.75 ;
END VIA12_4

VIA VIA23_1 DEFAULT
	LAYER METAL2 ;
		RECT -0.3 -0.3 0.3 0.3 ;
	LAYER VIA23 ;
		RECT -0.15 -0.15 0.15 0.15 ;
	LAYER METAL3 ;
		RECT -0.3 -0.3 0.3 0.3 ;
END VIA23_1

VIA VIA23_2H DEFAULT
	LAYER METAL2 ;
		RECT -0.75 -0.3 0.75 0.3 ;
	LAYER VIA23 ;
		RECT -0.6 -0.15 -0.3 0.15 ;
		RECT 0.3 -0.15 0.6 0.15 ;
	LAYER METAL3 ;
		RECT -0.75 -0.3 0.75 0.3 ;
END VIA23_2H

VIA VIA23_2V DEFAULT
	LAYER METAL2 ;
		RECT -0.3 -0.75 0.3 0.75 ;
	LAYER VIA23 ;
		RECT -0.15 -0.6 0.15 -0.3 ;
		RECT -0.15 0.3 0.15 0.6 ;
	LAYER METAL3 ;
		RECT -0.3 -0.75 0.3 0.75 ;
END VIA23_2V

VIA VIA23_4 DEFAULT
	LAYER METAL2 ;
		RECT -0.75 -0.75 0.75 0.75 ;
	LAYER VIA23 ;
		RECT -0.6 -0.6 -0.3 -0.3 ;
		RECT -0.6 0.3 -0.3 0.6 ;
		RECT 0.3 0.3 0.6 0.6 ;
		RECT 0.3 -0.6 0.6 -0.3 ;
	LAYER METAL3 ;
		RECT -0.75 -0.75 0.75 0.75 ;
END VIA23_4

VIA VIA34_1 DEFAULT
	LAYER METAL3 ;
		RECT -0.3 -0.3 0.3 0.3 ;
	LAYER VIA34 ;
		RECT -0.15 -0.15 0.15 0.15 ;
	LAYER METAL4 ;
		RECT -0.3 -0.3 0.3 0.3 ;
END VIA34_1

VIA VIA34_2H DEFAULT
	LAYER METAL3 ;
		RECT -0.75 -0.3 0.75 0.3 ;
	LAYER VIA34 ;
		RECT -0.6 -0.15 -0.3 0.15 ;
		RECT 0.3 -0.15 0.6 0.15 ;
	LAYER METAL4 ;
		RECT -0.75 -0.3 0.75 0.3 ;
END VIA34_2H

VIA VIA34_2V DEFAULT
	LAYER METAL3 ;
		RECT -0.3 -0.75 0.3 0.75 ;
	LAYER VIA34 ;
		RECT -0.15 -0.6 0.15 -0.3 ;
		RECT -0.15 0.3 0.15 0.6 ;
	LAYER METAL4 ;
		RECT -0.3 -0.75 0.3 0.75 ;
END VIA34_2V

VIA VIA34_4 DEFAULT
	LAYER METAL3 ;
		RECT -0.75 -0.75 0.75 0.75 ;
	LAYER VIA34 ;
		RECT -0.6 -0.6 -0.3 -0.3 ;
		RECT -0.6 0.3 -0.3 0.6 ;
		RECT 0.3 0.3 0.6 0.6 ;
		RECT 0.3 -0.6 0.6 -0.3 ;
	LAYER METAL4 ;
		RECT -0.75 -0.75 0.75 0.75 ;
END VIA34_4

VIA VIA45_1 DEFAULT
	LAYER METAL4 ;
		RECT -1.8 -1.8 1.8 1.8 ;
	LAYER VIA45 ;
		RECT -1.2 -1.2 1.2 1.2 ;
	LAYER RDL ;
		RECT -1.8 -1.8 1.8 1.8 ;
END VIA45_1

VIARULE VIA_GEN_12 GENERATE
	LAYER METAL1 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER METAL2 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER VIA12 ;
	RECT -0.15 -0.15 0.15 0.15 ;
	SPACING 0.6 BY 0.6 ;
END VIA_GEN_12

VIARULE VIA_GEN_23 GENERATE
	LAYER METAL2 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER METAL3 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER VIA23 ;
	RECT -0.15 -0.15 0.15 0.15 ;
	SPACING 0.6 BY 0.6 ;
END VIA_GEN_23

VIARULE VIA_GEN_34 GENERATE
	LAYER METAL3 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER METAL4 ;
	ENCLOSURE 0.15 0.15 ;
	WIDTH 0.3 TO 15 ;
	LAYER VIA34 ;
	RECT -0.15 -0.15 0.15 0.15 ;
	SPACING 0.6 BY 0.6 ;
END VIA_GEN_34

VIARULE VIA_GEN_45 GENERATE
	LAYER METAL4 ;
	ENCLOSURE 0.6 0.6 ;
	WIDTH 0.3 TO 15 ;
	LAYER RDL ;
	ENCLOSURE 0.6 0.6 ;
	WIDTH 2.8 TO 30.0 ;
	LAYER VIA45 ;
	RECT -1.2 -1.2 1.2 1.2 ;
	SPACING 4.8 BY 4.8 ;
END VIA_GEN_45

SITE CORE0
	SIZE 0.3 BY 1.5 ;
	CLASS CORE ;
	SYMMETRY X Y  ;
END CORE0

