VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO UBUMP
	CLASS COVER BUMP ;
	ORIGIN 0 0 ;
	SIZE 22.5 BY 22.5 ;
	SYMMETRY X Y ;
	PIN PAD
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER RDL ;
				POLYGON 6.59 0 15.91 0 22.5 6.59 22.5 15.91 15.91 22.5 6.59 22.5 0 15.91 0 6.59 ; 
		END
	END PAD
	OBS
		LAYER VIA45 SPACING 0.000 ;
			POLYGON 6.59 2 15.91 2 20.5 6.59 20.5 15.91 15.91 20.5 6.59 20.5 2 15.91 2 6.59 ; 
	END
END UBUMP

MACRO C4BUMP
	CLASS COVER BUMP ;
	ORIGIN 0 0 ;
	SIZE 70 BY 70 ;
	SYMMETRY X Y ;
	PIN PAD
		DIRECTION INOUT ;
		USE SIGNAL ;
		PORT
			LAYER MB ;
		    		POLYGON 20.5025 0 49.4975 0 70 20.5025 70 49.4975 49.4975 70 20.5025 70 0 49.4975 0 20.5025 ;
		  	LAYER TSV1 ;
		    		RECT 25 23 45 47 ;
		  	LAYER METAL1 ;
		    		RECT 22 20 48 50 ;
		END
	END PAD
	OBS
	  	LAYER METAL1 SPACING 0.000 ;
	    		RECT 20 18 50 19 ;
	    		RECT 20 51 50 52 ;
	    		RECT 20 18 21 51 ;
	    		RECT 49 18 50 51 ;
	END
END C4BUMP

END LIBRARY

